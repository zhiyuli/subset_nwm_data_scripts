netcdf nwm.t00z.analysis_assim.terrain_rt.tm00.conus {
dimensions:
	time = UNLIMITED ; // (1 currently)
	x = 18432 ;
	y = 15360 ;
	reference_time = 1 ;
variables:
	int time(time) ;
		time:long_name = "valid output time" ;
		time:standard_name = "time" ;
		time:units = "minutes since 1970-01-01 00:00:00 UTC" ;
		time:_Storage = "chunked" ;
		time:_ChunkSizes = 1048576 ;
		time:_DeflateLevel = 2 ;
		time:_Shuffle = "true" ;
		time:_Endianness = "little" ;
	int zwattablrt(time, y, x) ;
		zwattablrt:_FillValue = -99990 ;
		zwattablrt:units = "m" ;
		zwattablrt:long_name = "water table depth" ;
		zwattablrt:grid_mapping = "ProjectionCoordinateSystem" ;
		zwattablrt:proj4 = "+proj=lcc +lat_1=30 +lat_2=60 +lat_0=40 +lon_0=-97 +x_0=0 +y_0=0 +a=6370000 +b=6370000 +units=m +no_defs" ;
		zwattablrt:esri_pe_string = "PROJCS[\"Sphere_Lambert_Conformal_Conic\",GEOGCS[\"GCS_Sphere\",DATUM[\"D_Sphere\",SPHEROID[\"Sphere\",6370000.0,0.0]],PRIMEM[\"Greenwich\",0.0],UNIT[\"Degree\",0.0174532925199433]],PROJECTION[\"Lambert_Conformal_Conic\"],PARAMETER[\"false_easting\",0.0],PARAMETER[\"false_northing\",0.0],PARAMETER[\"central_meridian\",-97.0],PARAMETER[\"standard_parallel_1\",30.0],PARAMETER[\"standard_parallel_2\",60.0],PARAMETER[\"latitude_of_origin\",40.0000076294],UNIT[\"Meter\",1.0]];-35691800 -29075200 126180232.640845;-100000 10000;-100000 10000;0.001;0.001;0.001;IsHighPrecision" ;
		zwattablrt:scale_factor = 0.1 ;
		zwattablrt:add_offset = 0. ;
		zwattablrt:valid_range = 0., 100. ;
		zwattablrt:missing_value = -99990 ;
		zwattablrt:_Storage = "chunked" ;
		zwattablrt:_ChunkSizes = 1, 904, 1085 ;
		zwattablrt:_DeflateLevel = 2 ;
		zwattablrt:_Shuffle = "true" ;
		zwattablrt:_Endianness = "little" ;
	int sfcheadsubrt(time, y, x) ;
		sfcheadsubrt:_FillValue = -9999 ;
		sfcheadsubrt:units = "mm" ;
		sfcheadsubrt:long_name = "surface head" ;
		sfcheadsubrt:grid_mapping = "ProjectionCoordinateSystem" ;
		sfcheadsubrt:proj4 = "+proj=lcc +lat_1=30 +lat_2=60 +lat_0=40 +lon_0=-97 +x_0=0 +y_0=0 +a=6370000 +b=6370000 +units=m +no_defs" ;
		sfcheadsubrt:esri_pe_string = "PROJCS[\"Sphere_Lambert_Conformal_Conic\",GEOGCS[\"GCS_Sphere\",DATUM[\"D_Sphere\",SPHEROID[\"Sphere\",6370000.0,0.0]],PRIMEM[\"Greenwich\",0.0],UNIT[\"Degree\",0.0174532925199433]],PROJECTION[\"Lambert_Conformal_Conic\"],PARAMETER[\"false_easting\",0.0],PARAMETER[\"false_northing\",0.0],PARAMETER[\"central_meridian\",-97.0],PARAMETER[\"standard_parallel_1\",30.0],PARAMETER[\"standard_parallel_2\",60.0],PARAMETER[\"latitude_of_origin\",40.0000076294],UNIT[\"Meter\",1.0]];-35691800 -29075200 126180232.640845;-100000 10000;-100000 10000;0.001;0.001;0.001;IsHighPrecision" ;
		sfcheadsubrt:scale_factor = 1. ;
		sfcheadsubrt:add_offset = 0. ;
		sfcheadsubrt:valid_range = 0., 1000000. ;
		sfcheadsubrt:missing_value = -9999 ;
		sfcheadsubrt:_Storage = "chunked" ;
		sfcheadsubrt:_ChunkSizes = 1, 904, 1085 ;
		sfcheadsubrt:_DeflateLevel = 2 ;
		sfcheadsubrt:_Shuffle = "true" ;
		sfcheadsubrt:_Endianness = "little" ;
	int x_index(y, x) ;
		x_index:_FillValue = -9999 ;
		x_index:units = "mm" ;
		x_index:long_name = "x_index" ;
		x_index:grid_mapping = "ProjectionCoordinateSystem" ;
		x_index:proj4 = "+proj=lcc +lat_1=30 +lat_2=60 +lat_0=40 +lon_0=-97 +x_0=0 +y_0=0 +a=6370000 +b=6370000 +units=m +no_defs" ;
		x_index:esri_pe_string = "PROJCS[\"Sphere_Lambert_Conformal_Conic\",GEOGCS[\"GCS_Sphere\",DATUM[\"D_Sphere\",SPHEROID[\"Sphere\",6370000.0,0.0]],PRIMEM[\"Greenwich\",0.0],UNIT[\"Degree\",0.0174532925199433]],PROJECTION[\"Lambert_Conformal_Conic\"],PARAMETER[\"false_easting\",0.0],PARAMETER[\"false_northing\",0.0],PARAMETER[\"central_meridian\",-97.0],PARAMETER[\"standard_parallel_1\",30.0],PARAMETER[\"standard_parallel_2\",60.0],PARAMETER[\"latitude_of_origin\",40.0000076294],UNIT[\"Meter\",1.0]];-35691800 -29075200 126180232.640845;-100000 10000;-100000 10000;0.001;0.001;0.001;IsHighPrecision" ;		
		x_index:_Storage = "chunked" ;
		x_index:_ChunkSizes = 904, 1085 ;
		x_index:_DeflateLevel = 2 ;
		x_index:_Shuffle = "true" ;
		x_index:_Endianness = "little" ;
	int y_index(y, x) ;
		y_index:_FillValue = -9999 ;
		y_index:units = "mm" ;
		y_index:long_name = "y_index" ;
		y_index:grid_mapping = "ProjectionCoordinateSystem" ;
		y_index:proj4 = "+proj=lcc +lat_1=30 +lat_2=60 +lat_0=40 +lon_0=-97 +x_0=0 +y_0=0 +a=6370000 +b=6370000 +units=m +no_defs" ;
		y_index:esri_pe_string = "PROJCS[\"Sphere_Lambert_Conformal_Conic\",GEOGCS[\"GCS_Sphere\",DATUM[\"D_Sphere\",SPHEROID[\"Sphere\",6370000.0,0.0]],PRIMEM[\"Greenwich\",0.0],UNIT[\"Degree\",0.0174532925199433]],PROJECTION[\"Lambert_Conformal_Conic\"],PARAMETER[\"false_easting\",0.0],PARAMETER[\"false_northing\",0.0],PARAMETER[\"central_meridian\",-97.0],PARAMETER[\"standard_parallel_1\",30.0],PARAMETER[\"standard_parallel_2\",60.0],PARAMETER[\"latitude_of_origin\",40.0000076294],UNIT[\"Meter\",1.0]];-35691800 -29075200 126180232.640845;-100000 10000;-100000 10000;0.001;0.001;0.001;IsHighPrecision" ;		
		y_index:_Storage = "chunked" ;
		y_index:_ChunkSizes = 904, 1085 ;
		y_index:_DeflateLevel = 2 ;
		y_index:_Shuffle = "true" ;
		y_index:_Endianness = "little" ;
	double x(x) ;
		x:standard_name = "projection_x_coordinate" ;
		x:long_name = "x coordinate of projection" ;
		x:_CoordinateAxisType = "GeoX" ;
		x:units = "m" ;
		x:resolution = 250. ;
		x:_Storage = "chunked" ;
		x:_ChunkSizes = 18432 ;
		x:_DeflateLevel = 2 ;
		x:_Shuffle = "true" ;
		x:_Endianness = "little" ;	
	double y(y) ;
		y:standard_name = "projection_y_coordinate" ;
		y:long_name = "y coordinate of projection" ;
		y:_CoordinateAxisType = "GeoY" ;
		y:units = "m" ;
		y:resolution = 250. ;
		y:_Storage = "chunked" ;
		y:_ChunkSizes = 15360 ;
		y:_DeflateLevel = 2 ;
		y:_Shuffle = "true" ;
		y:_Endianness = "little" ;	
	char ProjectionCoordinateSystem ;
		ProjectionCoordinateSystem:_CoordinateTransformType = "Projection" ;
		ProjectionCoordinateSystem:transform_name = "lambert_conformal_conic" ;
		ProjectionCoordinateSystem:grid_mapping_name = "lambert_conformal_conic" ;
		ProjectionCoordinateSystem:_CoordinateAxes = "y x" ;
		ProjectionCoordinateSystem:esri_pe_string = "PROJCS[\"Sphere_Lambert_Conformal_Conic\",GEOGCS[\"GCS_Sphere\",DATUM[\"D_Sphere\",SPHEROID[\"Sphere\",6370000.0,0.0]],PRIMEM[\"Greenwich\",0.0],UNIT[\"Degree\",0.0174532925199433]],PROJECTION[\"Lambert_Conformal_Conic\"],PARAMETER[\"false_easting\",0.0],PARAMETER[\"false_northing\",0.0],PARAMETER[\"central_meridian\",-97.0],PARAMETER[\"standard_parallel_1\",30.0],PARAMETER[\"standard_parallel_2\",60.0],PARAMETER[\"latitude_of_origin\",40.0000076294],UNIT[\"Meter\",1.0]];-35691800 -29075200 126180232.640845;-100000 10000;-100000 10000;0.001;0.001;0.001;IsHighPrecision" ;
		ProjectionCoordinateSystem:standard_parallel = 30., 60. ;
		ProjectionCoordinateSystem:longitude_of_central_meridian = -97. ;
		ProjectionCoordinateSystem:latitude_of_projection_origin = 40.0000076294 ;
		ProjectionCoordinateSystem:false_easting = 0. ;
		ProjectionCoordinateSystem:false_northing = 0. ;
		ProjectionCoordinateSystem:earth_radius = 6370000. ;
		ProjectionCoordinateSystem:proj4 = "+proj=lcc +lat_1=30 +lat_2=60 +lat_0=40 +lon_0=-97 +x_0=0 +y_0=0 +a=6370000 +b=6370000 +units=m +no_defs" ;
	int reference_time(reference_time) ;
		reference_time:long_name = "model initialization time" ;
		reference_time:standard_name = "forecast_reference_time" ;
		reference_time:units = "minutes since 1970-01-01 00:00:00 UTC" ;
		reference_time:_Storage = "contiguous" ;
		reference_time:_Endianness = "little" ;

// global attributes:
		:model_initialization_time = "2017-04-01_21:00:00" ;
		:model_output_valid_time = "2017-04-02_00:00:00" ;
		:output_decimation_factor = 1 ;
		:Conventions = "CF-1.6" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4 classic model" ;
}
